entity Testbench is 
end Testbench;

architecture tb of Testbench is
	signal s_0,s_1,a_0,a_1,a_2,a_3,a_4,a_5,a_6,a_7,a_8,a_9,a_10,a_11,a_12,a_13,a_14,a_15,
	b_0,b_1,b_2,b_3,b_4,b_5,b_6,b_7,b_8,b_9,b_10,b_11,b_12,b_13,b_14,b_15 : bit;
	signal c_0,c_1,c_2,c_3,c_4,c_5,c_6,c_7,c_8,c_9,c_10,c_11,c_12,c_13,c_14,c_15,c_,z_: bit;
	
	component ALU is 
		port(S0,S1,A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15, B0, B1, B2, B3, B4, B5, B6, B7, B8, B9, B10, B11, B12, B13, B14, B15: in bit;
			C0, C1, C2, C3, C4, C5, C6, C7, C8, C9, C10, C11, C12, C13, C14, C15,C,Z:out bit);
	end component;
	
	begin
	dut_instance: ALU
	port map(s_0,s_1,a_0,a_1,a_2,a_3,a_4,a_5,a_6,a_7,a_8,a_9,a_10,a_11,a_12,a_13,a_14,a_15,
	b_0,b_1,b_2,b_3,b_4,b_5,b_6,b_7,b_8,b_9,b_10,b_11,b_12,b_13,b_14,b_15,
	c_0,c_1,c_2,c_3,c_4,c_5,c_6,c_7,c_8,c_9,c_10,c_11,c_12,c_13,c_14,c_15,c_,z_);

	process
	begin
		
		s_0 <= '0';
		s_1 <= '0';
		a_0 <= '0';
		a_1 <= '0';
		a_2 <= '0';
		a_3 <= '0';
		a_4 <= '0';
		a_5 <= '0';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '0';
		a_11 <= '0';
		a_12 <= '0';
		a_13 <= '0';
		a_14 <= '0';
		a_15 <= '0';
		b_0 <= '0';
		b_1 <= '0';
		b_2 <= '0';
		b_3 <= '0';
		b_4 <= '0';
		b_5 <= '0';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '0';
		b_11 <= '0';
		b_12 <= '0';
		b_13 <= '0';
		b_14 <= '0';
		b_15 <= '0';
		
		wait for 10 ns;
		
		s_0 <= '0';
		s_1 <= '0';
		a_0 <= '1';
		a_1 <= '1';
		a_2 <= '1';
		a_3 <= '1';
		a_4 <= '1';
		a_5 <= '1';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '0';
		a_11 <= '0';
		a_12 <= '0';
		a_13 <= '0';
		a_14 <= '0';
		a_15 <= '0';
		b_0 <= '0';
		b_1 <= '0';
		b_2 <= '0';
		b_3 <= '0';
		b_4 <= '0';
		b_5 <= '0';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '0';
		b_11 <= '0';
		b_12 <= '0';
		b_13 <= '0';
		b_14 <= '0';
		b_15 <= '0';
		
		wait for 10 ns;
		
		s_0 <= '0';
		s_1 <= '0';
		a_0 <= '1'
a_1 <= '1';
a_2 <= '1';
a_3 <= '1';
a_4 <= '1';
a_5 <= '1';
a_6 <= '1';
a_7 <= '1';
a_8 <= '1';
a_9 <= '1';
a_10 <= '1';
a_11 <= '1';
a_12 <= '1';
a_13 <= '1';
a_14 <= '1';
a_15 <= '1';
b_0 <= '1';
b_1 <= '1';
b_2 <= '1';
b_3 <= '1';
b_4 <= '1';
b_5 <= '1';
b_6 <= '1';
b_7 <= '1';
b_8 <= '1';
b_9 <= '1';
b_10 <= '1';
b_11 <= '1';
b_12 <= '1';
b_13 <= '1';
b_14 <= '1';
b_15 <= '1';

wait for 10 ns;

s_0 <= '0';
		s_1 <= '0';
		a_0 <= '0';
		a_1 <= '0';
		a_2 <= '0';
		a_3 <= '0';
		a_4 <= '0';
		a_5 <= '0';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '0';
		a_11 <= '0';
		a_12 <= '0';
		a_13 <= '0';
		a_14 <= '0';
		a_15 <= '0';
		b_0 <= '1';
		b_1 <= '1';
		b_2 <= '1';
		b_3 <= '1';
		b_4 <= '1';
		b_5 <= '1';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '0';
		b_11 <= '0';
		b_12 <= '0';
		b_13 <= '0';
		b_14 <= '0';
		b_15 <= '0';
		
		wait for 10 ns;
		
		s_0 <= '0';
		s_1 <= '0';
		a_0 <= '0';
		a_1 <= '0';
		a_2 <= '0';
		a_3 <= '0';
		a_4 <= '0';
		a_5 <= '0';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '1';
		a_11 <= '1';
		a_12 <= '1';
		a_13 <= '1';
		a_14 <= '1';
		a_15 <= '1';
		b_0 <= '0';
		b_1 <= '0';
		b_2 <= '0';
		b_3 <= '0';
		b_4 <= '0';
		b_5 <= '0';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '1';
		b_11 <= '1';
		b_12 <= '1';
		b_13 <= '1';
		b_14 <= '1';
		b_15 <= '1';
		
		wait for 10 ns;
		
		s_0 <= '0';
		s_1 <= '1';
		a_0 <= '0';
		a_1 <= '0';
		a_2 <= '0';
		a_3 <= '0';
		a_4 <= '0';
		a_5 <= '0';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '0';
		a_11 <= '0';
		a_12 <= '0';
		a_13 <= '0';
		a_14 <= '0';
		a_15 <= '0';
		b_0 <= '0';
		b_1 <= '0';
		b_2 <= '0';
		b_3 <= '0';
		b_4 <= '0';
		b_5 <= '0';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '0';
		b_11 <= '0';
		b_12 <= '0';
		b_13 <= '0';
		b_14 <= '0';
		b_15 <= '0';
		
		wait for 10 ns;
		
		s_0 <= '0';
		s_1 <= '1';
		a_0 <= '1';
		a_1 <= '1';
		a_2 <= '1';
		a_3 <= '1';
		a_4 <= '1';
		a_5 <= '1';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '0';
		a_11 <= '0';
		a_12 <= '0';
		a_13 <= '0';
		a_14 <= '0';
		a_15 <= '0';
		b_0 <= '0';
		b_1 <= '0';
		b_2 <= '0';
		b_3 <= '0';
		b_4 <= '0';
		b_5 <= '0';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '0';
		b_11 <= '0';
		b_12 <= '0';
		b_13 <= '0';
		b_14 <= '0';
		b_15 <= '0';
		
		wait for 10 ns;
		
		s_0 <= '0';
		s_1 <= '1';
		a_0 <= '1'
a_1 <= '1';
a_2 <= '1';
a_3 <= '1';
a_4 <= '1';
a_5 <= '1';
a_6 <= '1';
a_7 <= '1';
a_8 <= '1';
a_9 <= '1';
a_10 <= '1';
a_11 <= '1';
a_12 <= '1';
a_13 <= '1';
a_14 <= '1';
a_15 <= '1';
b_0 <= '1';
b_1 <= '1';
b_2 <= '1';
b_3 <= '1';
b_4 <= '1';
b_5 <= '1';
b_6 <= '1';
b_7 <= '1';
b_8 <= '1';
b_9 <= '1';
b_10 <= '1';
b_11 <= '1';
b_12 <= '1';
b_13 <= '1';
b_14 <= '1';
b_15 <= '1';

wait for 10 ns;

		s_0 <= '0';
		s_1 <= '1';
		a_0 <= '0';
		a_1 <= '0';
		a_2 <= '0';
		a_3 <= '0';
		a_4 <= '0';
		a_5 <= '0';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '0';
		a_11 <= '0';
		a_12 <= '0';
		a_13 <= '0';
		a_14 <= '0';
		a_15 <= '0';
		b_0 <= '1';
		b_1 <= '1';
		b_2 <= '1';
		b_3 <= '1';
		b_4 <= '1';
		b_5 <= '1';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '0';
		b_11 <= '0';
		b_12 <= '0';
		b_13 <= '0';
		b_14 <= '0';
		b_15 <= '0';
		
		wait for 10 ns;
		
		s_0 <= '0';
		s_1 <= '1';
		a_0 <= '0';
		a_1 <= '0';
		a_2 <= '0';
		a_3 <= '0';
		a_4 <= '0';
		a_5 <= '0';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '1';
		a_11 <= '1';
		a_12 <= '1';
		a_13 <= '1';
		a_14 <= '1';
		a_15 <= '1';
		b_0 <= '0';
		b_1 <= '0';
		b_2 <= '0';
		b_3 <= '0';
		b_4 <= '0';
		b_5 <= '0';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '1';
		b_11 <= '1';
		b_12 <= '1';
		b_13 <= '1';
		b_14 <= '1';
		b_15 <= '1';
		
		wait for 10 ns;
		
		s_0 <= '1';
		s_1 <= '0';
		a_0 <= '0';
		a_1 <= '0';
		a_2 <= '0';
		a_3 <= '0';
		a_4 <= '0';
		a_5 <= '0';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '0';
		a_11 <= '0';
		a_12 <= '0';
		a_13 <= '0';
		a_14 <= '0';
		a_15 <= '0';
		b_0 <= '0';
		b_1 <= '0';
		b_2 <= '0';
		b_3 <= '0';
		b_4 <= '0';
		b_5 <= '0';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '0';
		b_11 <= '0';
		b_12 <= '0';
		b_13 <= '0';
		b_14 <= '0';
		b_15 <= '0';
		
		wait for 10 ns;
		
		s_0 <= '1';
		s_1 <= '0';
		a_0 <= '1';
		a_1 <= '1';
		a_2 <= '1';
		a_3 <= '1';
		a_4 <= '1';
		a_5 <= '1';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '0';
		a_11 <= '0';
		a_12 <= '0';
		a_13 <= '0';
		a_14 <= '0';
		a_15 <= '0';
		b_0 <= '0';
		b_1 <= '0';
		b_2 <= '0';
		b_3 <= '0';
		b_4 <= '0';
		b_5 <= '0';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '0';
		b_11 <= '0';
		b_12 <= '0';
		b_13 <= '0';
		b_14 <= '0';
		b_15 <= '0';
		
		wait for 10 ns;
		
		s_0 <= '1';
		s_1 <= '0';
		a_0 <= '1'
a_1 <= '1';
a_2 <= '1';
a_3 <= '1';
a_4 <= '1';
a_5 <= '1';
a_6 <= '1';
a_7 <= '1';
a_8 <= '1';
a_9 <= '1';
a_10 <= '1';
a_11 <= '1';
a_12 <= '1';
a_13 <= '1';
a_14 <= '1';
a_15 <= '1';
b_0 <= '1';
b_1 <= '1';
b_2 <= '1';
b_3 <= '1';
b_4 <= '1';
b_5 <= '1';
b_6 <= '1';
b_7 <= '1';
b_8 <= '1';
b_9 <= '1';
b_10 <= '1';
b_11 <= '1';
b_12 <= '1';
b_13 <= '1';
b_14 <= '1';
b_15 <= '1';

wait for 10 ns;

		s_0 <= '1';
		s_1 <= '0';
		a_0 <= '0';
		a_1 <= '0';
		a_2 <= '0';
		a_3 <= '0';
		a_4 <= '0';
		a_5 <= '0';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '0';
		a_11 <= '0';
		a_12 <= '0';
		a_13 <= '0';
		a_14 <= '0';
		a_15 <= '0';
		b_0 <= '1';
		b_1 <= '1';
		b_2 <= '1';
		b_3 <= '1';
		b_4 <= '1';
		b_5 <= '1';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '0';
		b_11 <= '0';
		b_12 <= '0';
		b_13 <= '0';
		b_14 <= '0';
		b_15 <= '0';
		
		wait for 10 ns;
		
		s_0 <= '1';
		s_1 <= '0';
		a_0 <= '0';
		a_1 <= '0';
		a_2 <= '0';
		a_3 <= '0';
		a_4 <= '0';
		a_5 <= '0';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '1';
		a_11 <= '1';
		a_12 <= '1';
		a_13 <= '1';
		a_14 <= '1';
		a_15 <= '1';
		b_0 <= '0';
		b_1 <= '0';
		b_2 <= '0';
		b_3 <= '0';
		b_4 <= '0';
		b_5 <= '0';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '1';
		b_11 <= '1';
		b_12 <= '1';
		b_13 <= '1';
		b_14 <= '1';
		b_15 <= '1';
		
		wait for 10 ns;
		
		s_0 <= '1';
		s_1 <= '1';
		a_0 <= '0';
		a_1 <= '0';
		a_2 <= '0';
		a_3 <= '0';
		a_4 <= '0';
		a_5 <= '0';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '0';
		a_11 <= '0';
		a_12 <= '0';
		a_13 <= '0';
		a_14 <= '0';
		a_15 <= '0';
		b_0 <= '0';
		b_1 <= '0';
		b_2 <= '0';
		b_3 <= '0';
		b_4 <= '0';
		b_5 <= '0';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '0';
		b_11 <= '0';
		b_12 <= '0';
		b_13 <= '0';
		b_14 <= '0';
		b_15 <= '0';
		
		wait for 10 ns;
		
		s_0 <= '1';
		s_1 <= '1';
		a_0 <= '1';
		a_1 <= '1';
		a_2 <= '1';
		a_3 <= '1';
		a_4 <= '1';
		a_5 <= '1';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '0';
		a_11 <= '0';
		a_12 <= '0';
		a_13 <= '0';
		a_14 <= '0';
		a_15 <= '0';
		b_0 <= '0';
		b_1 <= '0';
		b_2 <= '0';
		b_3 <= '0';
		b_4 <= '0';
		b_5 <= '0';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '0';
		b_11 <= '0';
		b_12 <= '0';
		b_13 <= '0';
		b_14 <= '0';
		b_15 <= '0';
		
		wait for 10 ns;
		
		s_0 <= '1';
		s_1 <= '1';
		a_0 <= '1'
a_1 <= '1';
a_2 <= '1';
a_3 <= '1';
a_4 <= '1';
a_5 <= '1';
a_6 <= '1';
a_7 <= '1';
a_8 <= '1';
a_9 <= '1';
a_10 <= '1';
a_11 <= '1';
a_12 <= '1';
a_13 <= '1';
a_14 <= '1';
a_15 <= '1';
b_0 <= '1';
b_1 <= '1';
b_2 <= '1';
b_3 <= '1';
b_4 <= '1';
b_5 <= '1';
b_6 <= '1';
b_7 <= '1';
b_8 <= '1';
b_9 <= '1';
b_10 <= '1';
b_11 <= '1';
b_12 <= '1';
b_13 <= '1';
b_14 <= '1';
b_15 <= '1';

wait for 10 ns;

		s_0 <= '1';
		s_1 <= '1';
		a_0 <= '0';
		a_1 <= '0';
		a_2 <= '0';
		a_3 <= '0';
		a_4 <= '0';
		a_5 <= '0';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '0';
		a_11 <= '0';
		a_12 <= '0';
		a_13 <= '0';
		a_14 <= '0';
		a_15 <= '0';
		b_0 <= '1';
		b_1 <= '1';
		b_2 <= '1';
		b_3 <= '1';
		b_4 <= '1';
		b_5 <= '1';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '0';
		b_11 <= '0';
		b_12 <= '0';
		b_13 <= '0';
		b_14 <= '0';
		b_15 <= '0';
		
		wait for 10 ns;
		
		s_0 <= '1';
		s_1 <= '1';
		a_0 <= '0';
		a_1 <= '0';
		a_2 <= '0';
		a_3 <= '0';
		a_4 <= '0';
		a_5 <= '0';
		a_6 <= '0';
		a_7 <= '0';
		a_8 <= '0';
		a_9 <= '0';
		a_10 <= '1';
		a_11 <= '1';
		a_12 <= '1';
		a_13 <= '1';
		a_14 <= '1';
		a_15 <= '1';
		b_0 <= '0';
		b_1 <= '0';
		b_2 <= '0';
		b_3 <= '0';
		b_4 <= '0';
		b_5 <= '0';
		b_6 <= '0';
		b_7 <= '0';
		b_8 <= '0';
		b_9 <= '0';
		b_10 <= '1';
		b_11 <= '1';
		b_12 <= '1';
		b_13 <= '1';
		b_14 <= '1';
		b_15 <= '1';
		
		wait for 10 ns;
		
		end process;

end tb;
